--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   13:30:17 03/28/2016
-- Design Name:   
-- Module Name:   D:/Git/DIG_Assignment1/Projeckt/Komponenter/TeenthSec/TEST_teenthSec.vhd
-- Project Name:  TeenthSec
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: TeenthSec
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TEST_teenthSec IS
END TEST_teenthSec;
 
ARCHITECTURE behavior OF TEST_teenthSec IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT TeenthSec
    PORT(
         BCD : 	IN  std_logic_vector(3 downto 0);
         LED : 	OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal BCD : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal LED : std_logic_vector(7 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 

 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: TeenthSec PORT MAP (
          BCD => BCD,
          LED => LED
        );


 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		BCD <= "0001";
		wait for 100 ns;
      BCD <= "0010";
		wait for 100 ns;
		BCD <= "0011";
		wait for 100 ns;
		BCD <= "0100";
		wait for 100 ns;
		BCD <= "0101";
		wait for 100 ns;
		BCD <= "0110";
		wait for 100 ns;
		BCD <= "0111";

      -- insert stimulus here 

      wait;
   end process;

END;
